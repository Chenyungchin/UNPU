module DNN_Core (
    
);

// ============ module instantiatiion =============
// weight memory

// LBPE x 6

// AFL x 6
    
endmodule